module atan(input logic [8:0] y, x,
           output logic [2:0] dir);
  logic s;
  assign s = y[8] ^ x[8];
  always_comb begin
    dir = 2'd0;
    case(x)
    8'd0 : begin
      if(y > 8'd0) begin
        if(y > 8'd0) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd1 : begin
      if(y > 8'd0) begin
        if(y > 8'd2) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd2 : begin
      if(y > 8'd0) begin
        if(y > 8'd4) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd3 : begin
      if(y > 8'd1) begin
        if(y > 8'd7) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd4 : begin
      if(y > 8'd1) begin
        if(y > 8'd9) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd5 : begin
      if(y > 8'd2) begin
        if(y > 8'd12) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd6 : begin
      if(y > 8'd2) begin
        if(y > 8'd14) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd7 : begin
      if(y > 8'd2) begin
        if(y > 8'd16) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd8 : begin
      if(y > 8'd3) begin
        if(y > 8'd19) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd9 : begin
      if(y > 8'd3) begin
        if(y > 8'd21) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd10 : begin
      if(y > 8'd4) begin
        if(y > 8'd24) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd11 : begin
      if(y > 8'd4) begin
        if(y > 8'd26) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd12 : begin
      if(y > 8'd4) begin
        if(y > 8'd28) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd13 : begin
      if(y > 8'd5) begin
        if(y > 8'd31) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd14 : begin
      if(y > 8'd5) begin
        if(y > 8'd33) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd15 : begin
      if(y > 8'd6) begin
        if(y > 8'd36) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd16 : begin
      if(y > 8'd6) begin
        if(y > 8'd38) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd17 : begin
      if(y > 8'd7) begin
        if(y > 8'd41) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd18 : begin
      if(y > 8'd7) begin
        if(y > 8'd43) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd19 : begin
      if(y > 8'd7) begin
        if(y > 8'd45) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd20 : begin
      if(y > 8'd8) begin
        if(y > 8'd48) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd21 : begin
      if(y > 8'd8) begin
        if(y > 8'd50) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd22 : begin
      if(y > 8'd9) begin
        if(y > 8'd53) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd23 : begin
      if(y > 8'd9) begin
        if(y > 8'd55) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd24 : begin
      if(y > 8'd9) begin
        if(y > 8'd57) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd25 : begin
      if(y > 8'd10) begin
        if(y > 8'd60) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd26 : begin
      if(y > 8'd10) begin
        if(y > 8'd62) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd27 : begin
      if(y > 8'd11) begin
        if(y > 8'd65) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd28 : begin
      if(y > 8'd11) begin
        if(y > 8'd67) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd29 : begin
      if(y > 8'd12) begin
        if(y > 8'd70) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd30 : begin
      if(y > 8'd12) begin
        if(y > 8'd72) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd31 : begin
      if(y > 8'd12) begin
        if(y > 8'd74) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd32 : begin
      if(y > 8'd13) begin
        if(y > 8'd77) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd33 : begin
      if(y > 8'd13) begin
        if(y > 8'd79) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd34 : begin
      if(y > 8'd14) begin
        if(y > 8'd82) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd35 : begin
      if(y > 8'd14) begin
        if(y > 8'd84) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd36 : begin
      if(y > 8'd14) begin
        if(y > 8'd86) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd37 : begin
      if(y > 8'd15) begin
        if(y > 8'd89) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd38 : begin
      if(y > 8'd15) begin
        if(y > 8'd91) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd39 : begin
      if(y > 8'd16) begin
        if(y > 8'd94) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd40 : begin
      if(y > 8'd16) begin
        if(y > 8'd96) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd41 : begin
      if(y > 8'd16) begin
        if(y > 8'd98) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd42 : begin
      if(y > 8'd17) begin
        if(y > 8'd101) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd43 : begin
      if(y > 8'd17) begin
        if(y > 8'd103) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd44 : begin
      if(y > 8'd18) begin
        if(y > 8'd106) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd45 : begin
      if(y > 8'd18) begin
        if(y > 8'd108) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd46 : begin
      if(y > 8'd19) begin
        if(y > 8'd111) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd47 : begin
      if(y > 8'd19) begin
        if(y > 8'd113) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd48 : begin
      if(y > 8'd19) begin
        if(y > 8'd115) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd49 : begin
      if(y > 8'd20) begin
        if(y > 8'd118) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd50 : begin
      if(y > 8'd20) begin
        if(y > 8'd120) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd51 : begin
      if(y > 8'd21) begin
        if(y > 8'd123) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd52 : begin
      if(y > 8'd21) begin
        if(y > 8'd125) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd53 : begin
      if(y > 8'd21) begin
        if(y > 8'd127) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd54 : begin
      if(y > 8'd22) begin
        if(y > 8'd130) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd55 : begin
      if(y > 8'd22) begin
        if(y > 8'd132) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd56 : begin
      if(y > 8'd23) begin
        if(y > 8'd135) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd57 : begin
      if(y > 8'd23) begin
        if(y > 8'd137) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd58 : begin
      if(y > 8'd24) begin
        if(y > 8'd140) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd59 : begin
      if(y > 8'd24) begin
        if(y > 8'd142) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd60 : begin
      if(y > 8'd24) begin
        if(y > 8'd144) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd61 : begin
      if(y > 8'd25) begin
        if(y > 8'd147) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd62 : begin
      if(y > 8'd25) begin
        if(y > 8'd149) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd63 : begin
      if(y > 8'd26) begin
        if(y > 8'd152) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd64 : begin
      if(y > 8'd26) begin
        if(y > 8'd154) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd65 : begin
      if(y > 8'd26) begin
        if(y > 8'd156) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd66 : begin
      if(y > 8'd27) begin
        if(y > 8'd159) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd67 : begin
      if(y > 8'd27) begin
        if(y > 8'd161) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd68 : begin
      if(y > 8'd28) begin
        if(y > 8'd164) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd69 : begin
      if(y > 8'd28) begin
        if(y > 8'd166) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd70 : begin
      if(y > 8'd28) begin
        if(y > 8'd168) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd71 : begin
      if(y > 8'd29) begin
        if(y > 8'd171) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd72 : begin
      if(y > 8'd29) begin
        if(y > 8'd173) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd73 : begin
      if(y > 8'd30) begin
        if(y > 8'd176) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd74 : begin
      if(y > 8'd30) begin
        if(y > 8'd178) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd75 : begin
      if(y > 8'd31) begin
        if(y > 8'd181) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd76 : begin
      if(y > 8'd31) begin
        if(y > 8'd183) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd77 : begin
      if(y > 8'd31) begin
        if(y > 8'd185) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd78 : begin
      if(y > 8'd32) begin
        if(y > 8'd188) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd79 : begin
      if(y > 8'd32) begin
        if(y > 8'd190) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd80 : begin
      if(y > 8'd33) begin
        if(y > 8'd193) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd81 : begin
      if(y > 8'd33) begin
        if(y > 8'd195) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd82 : begin
      if(y > 8'd33) begin
        if(y > 8'd197) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd83 : begin
      if(y > 8'd34) begin
        if(y > 8'd200) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd84 : begin
      if(y > 8'd34) begin
        if(y > 8'd202) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd85 : begin
      if(y > 8'd35) begin
        if(y > 8'd205) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd86 : begin
      if(y > 8'd35) begin
        if(y > 8'd207) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd87 : begin
      if(y > 8'd36) begin
        if(y > 8'd210) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd88 : begin
      if(y > 8'd36) begin
        if(y > 8'd212) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd89 : begin
      if(y > 8'd36) begin
        if(y > 8'd214) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd90 : begin
      if(y > 8'd37) begin
        if(y > 8'd217) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd91 : begin
      if(y > 8'd37) begin
        if(y > 8'd219) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd92 : begin
      if(y > 8'd38) begin
        if(y > 8'd222) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd93 : begin
      if(y > 8'd38) begin
        if(y > 8'd224) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd94 : begin
      if(y > 8'd38) begin
        if(y > 8'd226) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd95 : begin
      if(y > 8'd39) begin
        if(y > 8'd229) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd96 : begin
      if(y > 8'd39) begin
        if(y > 8'd231) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd97 : begin
      if(y > 8'd40) begin
        if(y > 8'd234) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd98 : begin
      if(y > 8'd40) begin
        if(y > 8'd236) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd99 : begin
      if(y > 8'd41) begin
        if(y > 8'd239) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd100 : begin
      if(y > 8'd41) begin
        if(y > 8'd241) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd101 : begin
      if(y > 8'd41) begin
        if(y > 8'd243) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd102 : begin
      if(y > 8'd42) begin
        if(y > 8'd246) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd103 : begin
      if(y > 8'd42) begin
        if(y > 8'd248) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd104 : begin
      if(y > 8'd43) begin
        if(y > 8'd251) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd105 : begin
      if(y > 8'd43) begin
        if(y > 8'd253) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd106 : begin
      if(y > 8'd43) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd107 : begin
      if(y > 8'd44) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd108 : begin
      if(y > 8'd44) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd109 : begin
      if(y > 8'd45) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd110 : begin
      if(y > 8'd45) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd111 : begin
      if(y > 8'd45) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd112 : begin
      if(y > 8'd46) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd113 : begin
      if(y > 8'd46) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd114 : begin
      if(y > 8'd47) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd115 : begin
      if(y > 8'd47) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd116 : begin
      if(y > 8'd48) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd117 : begin
      if(y > 8'd48) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd118 : begin
      if(y > 8'd48) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd119 : begin
      if(y > 8'd49) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd120 : begin
      if(y > 8'd49) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd121 : begin
      if(y > 8'd50) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd122 : begin
      if(y > 8'd50) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd123 : begin
      if(y > 8'd50) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd124 : begin
      if(y > 8'd51) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd125 : begin
      if(y > 8'd51) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd126 : begin
      if(y > 8'd52) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd127 : begin
      if(y > 8'd52) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd128 : begin
      if(y > 8'd53) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd129 : begin
      if(y > 8'd53) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd130 : begin
      if(y > 8'd53) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd131 : begin
      if(y > 8'd54) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd132 : begin
      if(y > 8'd54) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd133 : begin
      if(y > 8'd55) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd134 : begin
      if(y > 8'd55) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd135 : begin
      if(y > 8'd55) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd136 : begin
      if(y > 8'd56) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd137 : begin
      if(y > 8'd56) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd138 : begin
      if(y > 8'd57) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd139 : begin
      if(y > 8'd57) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd140 : begin
      if(y > 8'd57) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd141 : begin
      if(y > 8'd58) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd142 : begin
      if(y > 8'd58) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd143 : begin
      if(y > 8'd59) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd144 : begin
      if(y > 8'd59) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd145 : begin
      if(y > 8'd60) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd146 : begin
      if(y > 8'd60) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd147 : begin
      if(y > 8'd60) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd148 : begin
      if(y > 8'd61) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd149 : begin
      if(y > 8'd61) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd150 : begin
      if(y > 8'd62) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd151 : begin
      if(y > 8'd62) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd152 : begin
      if(y > 8'd62) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd153 : begin
      if(y > 8'd63) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd154 : begin
      if(y > 8'd63) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd155 : begin
      if(y > 8'd64) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd156 : begin
      if(y > 8'd64) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd157 : begin
      if(y > 8'd65) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd158 : begin
      if(y > 8'd65) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd159 : begin
      if(y > 8'd65) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd160 : begin
      if(y > 8'd66) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd161 : begin
      if(y > 8'd66) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd162 : begin
      if(y > 8'd67) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd163 : begin
      if(y > 8'd67) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd164 : begin
      if(y > 8'd67) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd165 : begin
      if(y > 8'd68) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd166 : begin
      if(y > 8'd68) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd167 : begin
      if(y > 8'd69) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd168 : begin
      if(y > 8'd69) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd169 : begin
      if(y > 8'd70) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd170 : begin
      if(y > 8'd70) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd171 : begin
      if(y > 8'd70) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd172 : begin
      if(y > 8'd71) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd173 : begin
      if(y > 8'd71) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd174 : begin
      if(y > 8'd72) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd175 : begin
      if(y > 8'd72) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd176 : begin
      if(y > 8'd72) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd177 : begin
      if(y > 8'd73) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd178 : begin
      if(y > 8'd73) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd179 : begin
      if(y > 8'd74) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd180 : begin
      if(y > 8'd74) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd181 : begin
      if(y > 8'd74) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd182 : begin
      if(y > 8'd75) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd183 : begin
      if(y > 8'd75) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd184 : begin
      if(y > 8'd76) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd185 : begin
      if(y > 8'd76) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd186 : begin
      if(y > 8'd77) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd187 : begin
      if(y > 8'd77) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd188 : begin
      if(y > 8'd77) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd189 : begin
      if(y > 8'd78) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd190 : begin
      if(y > 8'd78) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd191 : begin
      if(y > 8'd79) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd192 : begin
      if(y > 8'd79) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd193 : begin
      if(y > 8'd79) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd194 : begin
      if(y > 8'd80) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd195 : begin
      if(y > 8'd80) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd196 : begin
      if(y > 8'd81) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd197 : begin
      if(y > 8'd81) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd198 : begin
      if(y > 8'd82) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd199 : begin
      if(y > 8'd82) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd200 : begin
      if(y > 8'd82) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd201 : begin
      if(y > 8'd83) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd202 : begin
      if(y > 8'd83) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd203 : begin
      if(y > 8'd84) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd204 : begin
      if(y > 8'd84) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd205 : begin
      if(y > 8'd84) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd206 : begin
      if(y > 8'd85) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd207 : begin
      if(y > 8'd85) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd208 : begin
      if(y > 8'd86) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd209 : begin
      if(y > 8'd86) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd210 : begin
      if(y > 8'd86) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd211 : begin
      if(y > 8'd87) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd212 : begin
      if(y > 8'd87) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd213 : begin
      if(y > 8'd88) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd214 : begin
      if(y > 8'd88) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd215 : begin
      if(y > 8'd89) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd216 : begin
      if(y > 8'd89) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd217 : begin
      if(y > 8'd89) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd218 : begin
      if(y > 8'd90) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd219 : begin
      if(y > 8'd90) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd220 : begin
      if(y > 8'd91) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd221 : begin
      if(y > 8'd91) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd222 : begin
      if(y > 8'd91) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd223 : begin
      if(y > 8'd92) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd224 : begin
      if(y > 8'd92) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd225 : begin
      if(y > 8'd93) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd226 : begin
      if(y > 8'd93) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd227 : begin
      if(y > 8'd94) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd228 : begin
      if(y > 8'd94) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd229 : begin
      if(y > 8'd94) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd230 : begin
      if(y > 8'd95) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd231 : begin
      if(y > 8'd95) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd232 : begin
      if(y > 8'd96) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd233 : begin
      if(y > 8'd96) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd234 : begin
      if(y > 8'd96) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd235 : begin
      if(y > 8'd97) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd236 : begin
      if(y > 8'd97) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd237 : begin
      if(y > 8'd98) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd238 : begin
      if(y > 8'd98) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd239 : begin
      if(y > 8'd98) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd240 : begin
      if(y > 8'd99) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd241 : begin
      if(y > 8'd99) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd242 : begin
      if(y > 8'd100) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd243 : begin
      if(y > 8'd100) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd244 : begin
      if(y > 8'd101) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd245 : begin
      if(y > 8'd101) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd246 : begin
      if(y > 8'd101) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd247 : begin
      if(y > 8'd102) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd248 : begin
      if(y > 8'd102) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd249 : begin
      if(y > 8'd103) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd250 : begin
      if(y > 8'd103) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd251 : begin
      if(y > 8'd103) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd252 : begin
      if(y > 8'd104) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd253 : begin
      if(y > 8'd104) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd254 : begin
      if(y > 8'd105) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    8'd255 : begin
      if(y > 8'd105) begin
        if(y > 8'd255) begin
          dir = 2'd2;
        end else begin
          dir = s ? 2'd3 : 2'd1;
        end
      end else begin
        dir = 2'd0;
      end
    end
    endcase
  end
endmodule : atan
